`include "Opcode.vh"

module mem_control (
    input [6:0] opcode,
    input [2:0] fnc,
    
    output [31:0] mask,
    output 
);

endmodule